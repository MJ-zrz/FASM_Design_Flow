`timescale 1ns/1ns
module Dadda#(
	parameter	InputWidth 		= 	18				,
	parameter 	OutputWidth 	= 	32
)
(
	input				[InputWidth-1 : 0]				sum0				,
	input				[InputWidth-1 : 0]				sum1				,
	input				[InputWidth-1 : 0]				sum2				,
	input				[InputWidth-1 : 0]				sum3				,
	input				[InputWidth-1 : 0]				sum4				,
	input				[InputWidth-1 : 0]				sum5				,
	input				[InputWidth-1 : 0]				sum6				,
	input				[InputWidth-1 : 0]				sum7				,
	

	output				[OutputWidth-1 : 0]						vector0							,
	output				[OutputWidth-1 : 0]						vector1							   //
);

	wire		[0:0]				sum_column0				;
	wire		[0:0]				sum_column1				;
	wire		[1:0]				sum_column2				;
	wire		[1:0]				sum_column3				;
	wire		[2:0]				sum_column4				;
	wire		[2:0]				sum_column5				;
	wire		[3:0]				sum_column6				;
	wire		[3:0]				sum_column7				;
	wire		[4:0]				sum_column8				;
	wire		[4:0]				sum_column9				;
	wire		[5:0]				sum_column10				;
	wire		[5:0]				sum_column11				;
	wire		[6:0]				sum_column12				;
	wire		[6:0]				sum_column13				;
	wire		[7:0]				sum_column14				;
	wire		[7:0]				sum_column15				;
	wire		[8:0]				sum_column16				;
	wire		[7:0]				sum_column17				;
	wire		[6:0]				sum_column18				;
	wire		[6:0]				sum_column19				;
	wire		[5:0]				sum_column20				;
	wire		[5:0]				sum_column21				;
	wire		[4:0]				sum_column22				;
	wire		[4:0]				sum_column23				;
	wire		[3:0]				sum_column24				;
	wire		[3:0]				sum_column25				;
	wire		[2:0]				sum_column26				;
	wire		[2:0]				sum_column27				;
	wire		[1:0]				sum_column28				;
	wire		[1:0]				sum_column29				;
	wire		[0:0]				sum_column30				;
	wire		[1:0]				sum_column31				;


		wire		sum_column4_3				;
	wire		sum_column5_3				;
	wire		sum_column5_4				;
	wire		sum_column6_4				;
	wire		sum_column6_5				;
	wire		sum_column6_6				;
	wire		sum_column7_4				;
	wire		sum_column7_5				;
	wire		sum_column7_6				;
	wire		sum_column7_7				;
	wire		sum_column8_5				;
	wire		sum_column8_6				;
	wire		sum_column8_7				;
	wire		sum_column8_8				;
	wire		sum_column8_9				;
	wire		sum_column9_5				;
	wire		sum_column9_6				;
	wire		sum_column9_7				;
	wire		sum_column9_8				;
	wire		sum_column9_9				;
	wire		sum_column9_10				;
	wire		sum_column10_6				;
	wire		sum_column10_7				;
	wire		sum_column10_8				;
	wire		sum_column10_9				;
	wire		sum_column10_10				;
	wire		sum_column10_11				;
	wire		sum_column10_12				;
	wire		sum_column11_6				;
	wire		sum_column11_7				;
	wire		sum_column11_8				;
	wire		sum_column11_9				;
	wire		sum_column11_10				;
	wire		sum_column11_11				;
	wire		sum_column11_12				;
	wire		sum_column11_13				;
	wire		sum_column12_7				;
	wire		sum_column12_8				;
	wire		sum_column12_9				;
	wire		sum_column12_10				;
	wire		sum_column12_11				;
	wire		sum_column12_12				;
	wire		sum_column12_13				;
	wire		sum_column12_14				;
	wire		sum_column12_15				;
	wire		sum_column13_7				;
	wire		sum_column13_8				;
	wire		sum_column13_9				;
	wire		sum_column13_10				;
	wire		sum_column13_11				;
	wire		sum_column13_12				;
	wire		sum_column13_13				;
	wire		sum_column13_14				;
	wire		sum_column13_15				;
	wire		sum_column13_16				;
	wire		sum_column14_8				;
	wire		sum_column14_9				;
	wire		sum_column14_10				;
	wire		sum_column14_11				;
	wire		sum_column14_12				;
	wire		sum_column14_13				;
	wire		sum_column14_14				;
	wire		sum_column14_15				;
	wire		sum_column14_16				;
	wire		sum_column14_17				;
	wire		sum_column14_18				;
	wire		sum_column15_8				;
	wire		sum_column15_9				;
	wire		sum_column15_10				;
	wire		sum_column15_11				;
	wire		sum_column15_12				;
	wire		sum_column15_13				;
	wire		sum_column15_14				;
	wire		sum_column15_15				;
	wire		sum_column15_16				;
	wire		sum_column15_17				;
	wire		sum_column15_18				;
	wire		sum_column15_19				;
	wire		sum_column16_9				;
	wire		sum_column16_10				;
	wire		sum_column16_11				;
	wire		sum_column16_12				;
	wire		sum_column16_13				;
	wire		sum_column16_14				;
	wire		sum_column16_15				;
	wire		sum_column16_16				;
	wire		sum_column16_17				;
	wire		sum_column16_18				;
	wire		sum_column16_19				;
	wire		sum_column16_20				;
	wire		sum_column16_21				;
	wire		sum_column17_8				;
	wire		sum_column17_9				;
	wire		sum_column17_10				;
	wire		sum_column17_11				;
	wire		sum_column17_12				;
	wire		sum_column17_13				;
	wire		sum_column17_14				;
	wire		sum_column17_15				;
	wire		sum_column17_16				;
	wire		sum_column17_17				;
	wire		sum_column17_18				;
	wire		sum_column17_19				;
	wire		sum_column17_20				;
	wire		sum_column17_21				;
	wire		sum_column18_7				;
	wire		sum_column18_8				;
	wire		sum_column18_9				;
	wire		sum_column18_10				;
	wire		sum_column18_11				;
	wire		sum_column18_12				;
	wire		sum_column18_13				;
	wire		sum_column18_14				;
	wire		sum_column18_15				;
	wire		sum_column18_16				;
	wire		sum_column18_17				;
	wire		sum_column18_18				;
	wire		sum_column18_19				;
	wire		sum_column19_7				;
	wire		sum_column19_8				;
	wire		sum_column19_9				;
	wire		sum_column19_10				;
	wire		sum_column19_11				;
	wire		sum_column19_12				;
	wire		sum_column19_13				;
	wire		sum_column19_14				;
	wire		sum_column19_15				;
	wire		sum_column19_16				;
	wire		sum_column19_17				;
	wire		sum_column19_18				;
	wire		sum_column20_6				;
	wire		sum_column20_7				;
	wire		sum_column20_8				;
	wire		sum_column20_9				;
	wire		sum_column20_10				;
	wire		sum_column20_11				;
	wire		sum_column20_12				;
	wire		sum_column20_13				;
	wire		sum_column20_14				;
	wire		sum_column20_15				;
	wire		sum_column20_16				;
	wire		sum_column21_6				;
	wire		sum_column21_7				;
	wire		sum_column21_8				;
	wire		sum_column21_9				;
	wire		sum_column21_10				;
	wire		sum_column21_11				;
	wire		sum_column21_12				;
	wire		sum_column21_13				;
	wire		sum_column21_14				;
	wire		sum_column21_15				;
	wire		sum_column22_5				;
	wire		sum_column22_6				;
	wire		sum_column22_7				;
	wire		sum_column22_8				;
	wire		sum_column22_9				;
	wire		sum_column22_10				;
	wire		sum_column22_11				;
	wire		sum_column22_12				;
	wire		sum_column22_13				;
	wire		sum_column23_5				;
	wire		sum_column23_6				;
	wire		sum_column23_7				;
	wire		sum_column23_8				;
	wire		sum_column23_9				;
	wire		sum_column23_10				;
	wire		sum_column23_11				;
	wire		sum_column23_12				;
	wire		sum_column24_4				;
	wire		sum_column24_5				;
	wire		sum_column24_6				;
	wire		sum_column24_7				;
	wire		sum_column24_8				;
	wire		sum_column24_9				;
	wire		sum_column24_10				;
	wire		sum_column25_4				;
	wire		sum_column25_5				;
	wire		sum_column25_6				;
	wire		sum_column25_7				;
	wire		sum_column25_8				;
	wire		sum_column25_9				;
	wire		sum_column26_3				;
	wire		sum_column26_4				;
	wire		sum_column26_5				;
	wire		sum_column26_6				;
	wire		sum_column26_7				;
	wire		sum_column27_3				;
	wire		sum_column27_4				;
	wire		sum_column27_5				;
	wire		sum_column27_6				;
	wire		sum_column28_2				;
	wire		sum_column28_3				;
	wire		sum_column28_4				;
	wire		sum_column29_2				;
	wire		sum_column29_3				;
	wire		sum_column30_1				;


	assign		sum_column0				=		{sum0[0]}				;
	assign		sum_column1				=		{sum0[1]}				;
	assign		sum_column2				=		{sum0[2], sum1[0]}				;
	assign		sum_column3				=		{sum0[3], sum1[1]}				;
	assign		sum_column4				=		{sum0[4], sum1[2], sum2[0]}				;
	assign		sum_column5				=		{sum0[5], sum1[3], sum2[1]}				;
	assign		sum_column6				=		{sum0[6], sum1[4], sum2[2], sum3[0]}				;
	assign		sum_column7				=		{sum0[7], sum1[5], sum2[3], sum3[1]}				;
	assign		sum_column8				=		{sum0[8], sum1[6], sum2[4], sum3[2], sum4[0]}				;
	assign		sum_column9				=		{sum0[9], sum1[7], sum2[5], sum3[3], sum4[1]}				;
	assign		sum_column10				=		{sum0[10], sum1[8], sum2[6], sum3[4], sum4[2], sum5[0]}				;
	assign		sum_column11				=		{sum0[11], sum1[9], sum2[7], sum3[5], sum4[3], sum5[1]}				;
	assign		sum_column12				=		{sum0[12], sum1[10], sum2[8], sum3[6], sum4[4], sum5[2], sum6[0]}				;
	assign		sum_column13				=		{sum0[13], sum1[11], sum2[9], sum3[7], sum4[5], sum5[3], sum6[1]}				;
	assign		sum_column14				=		{sum0[14], sum1[12], sum2[10], sum3[8], sum4[6], sum5[4], sum6[2], sum7[0]}				;
	assign		sum_column15				=		{sum0[15], sum1[13], sum2[11], sum3[9], sum4[7], sum5[5], sum6[3], sum7[1]}				;
	assign		sum_column16				=		{1'b1, sum0[16], sum1[14], sum2[12], sum3[10], sum4[8], sum5[6], sum6[4], sum7[2]}				;
	assign		sum_column17				=		{sum0[17], sum1[15], sum2[13], sum3[11], sum4[9], sum5[7], sum6[5], sum7[3]}				;
	assign		sum_column18				=		{sum1[16], sum2[14], sum3[12], sum4[10], sum5[8], sum6[6], sum7[4]}				;
	assign		sum_column19				=		{sum1[17], sum2[15], sum3[13], sum4[11], sum5[9], sum6[7], sum7[5]}				;
	assign		sum_column20				=		{sum2[16], sum3[14], sum4[12], sum5[10], sum6[8], sum7[6]}				;
	assign		sum_column21				=		{sum2[17], sum3[15], sum4[13], sum5[11], sum6[9], sum7[7]}				;
	assign		sum_column22				=		{sum3[16], sum4[14], sum5[12], sum6[10], sum7[8]}				;
	assign		sum_column23				=		{sum3[17], sum4[15], sum5[13], sum6[11], sum7[9]}				;
	assign		sum_column24				=		{sum4[16], sum5[14], sum6[12], sum7[10]}				;
	assign		sum_column25				=		{sum4[17], sum5[15], sum6[13], sum7[11]}				;
	assign		sum_column26				=		{sum5[16], sum6[14], sum7[12]}				;
	assign		sum_column27				=		{sum5[17], sum6[15], sum7[13]}				;
	assign		sum_column28				=		{sum6[16], sum7[14]}				;
	assign		sum_column29				=		{sum6[17], sum7[15]}				;
	assign		sum_column30				=		{sum7[16]}				;
	assign		sum_column31				=		{1'b1, sum7[17]}				;
	

	
    HA HA_inst_0(
        .A              (sum_column4[0])            ,
        .B              (sum_column4[1])            ,
        .sum            (sum_column4_3)            ,
        .carry          (sum_column5_3)               //           
    );   
    
    FA FA_inst_1(
        .A              (sum_column5[0])            ,
        .B              (sum_column5[1])            ,
        .Cin            (sum_column5[2])            ,
        .sum            (sum_column5_4)            ,
        .carry          (sum_column6_4)               //           
    );    
    
    FA FA_inst_2(
        .A              (sum_column6[0])            ,
        .B              (sum_column6[1])            ,
        .Cin            (sum_column6[2])            ,
        .sum            (sum_column6_5)            ,
        .carry          (sum_column7_4)               //           
    );    
    
    FA FA_inst_3(
        .A              (sum_column7[0])            ,
        .B              (sum_column7[1])            ,
        .Cin            (sum_column7[2])            ,
        .sum            (sum_column7_5)            ,
        .carry          (sum_column8_5)               //           
    );    
    
    FA FA_inst_4(
        .A              (sum_column8[0])            ,
        .B              (sum_column8[1])            ,
        .Cin            (sum_column8[2])            ,
        .sum            (sum_column8_6)            ,
        .carry          (sum_column9_5)               //           
    );    
    
    FA FA_inst_5(
        .A              (sum_column9[0])            ,
        .B              (sum_column9[1])            ,
        .Cin            (sum_column9[2])            ,
        .sum            (sum_column9_6)            ,
        .carry          (sum_column10_6)               //           
    );    
    
    FA FA_inst_6(
        .A              (sum_column10[0])            ,
        .B              (sum_column10[1])            ,
        .Cin            (sum_column10[2])            ,
        .sum            (sum_column10_7)            ,
        .carry          (sum_column11_6)               //           
    );    
    
    FA FA_inst_7(
        .A              (sum_column11[0])            ,
        .B              (sum_column11[1])            ,
        .Cin            (sum_column11[2])            ,
        .sum            (sum_column11_7)            ,
        .carry          (sum_column12_7)               //           
    );    
    
    FA FA_inst_8(
        .A              (sum_column12[0])            ,
        .B              (sum_column12[1])            ,
        .Cin            (sum_column12[2])            ,
        .sum            (sum_column12_8)            ,
        .carry          (sum_column13_7)               //           
    );    
    
    FA FA_inst_9(
        .A              (sum_column13[0])            ,
        .B              (sum_column13[1])            ,
        .Cin            (sum_column13[2])            ,
        .sum            (sum_column13_8)            ,
        .carry          (sum_column14_8)               //           
    );    
    
    FA FA_inst_10(
        .A              (sum_column14[0])            ,
        .B              (sum_column14[1])            ,
        .Cin            (sum_column14[2])            ,
        .sum            (sum_column14_9)            ,
        .carry          (sum_column15_8)               //           
    );    
    
    FA FA_inst_11(
        .A              (sum_column15[0])            ,
        .B              (sum_column15[1])            ,
        .Cin            (sum_column15[2])            ,
        .sum            (sum_column15_9)            ,
        .carry          (sum_column16_9)               //           
    );    
    
    FA FA_inst_12(
        .A              (sum_column16[0])            ,
        .B              (sum_column16[1])            ,
        .Cin            (sum_column16[2])            ,
        .sum            (sum_column16_10)            ,
        .carry          (sum_column17_8)               //           
    );    
    
    FA FA_inst_13(
        .A              (sum_column17[0])            ,
        .B              (sum_column17[1])            ,
        .Cin            (sum_column17[2])            ,
        .sum            (sum_column17_9)            ,
        .carry          (sum_column18_7)               //           
    );    
    
    FA FA_inst_14(
        .A              (sum_column18[0])            ,
        .B              (sum_column18[1])            ,
        .Cin            (sum_column18[2])            ,
        .sum            (sum_column18_8)            ,
        .carry          (sum_column19_7)               //           
    );    
    
    FA FA_inst_15(
        .A              (sum_column19[0])            ,
        .B              (sum_column19[1])            ,
        .Cin            (sum_column19[2])            ,
        .sum            (sum_column19_8)            ,
        .carry          (sum_column20_6)               //           
    );    
    
    FA FA_inst_16(
        .A              (sum_column20[0])            ,
        .B              (sum_column20[1])            ,
        .Cin            (sum_column20[2])            ,
        .sum            (sum_column20_7)            ,
        .carry          (sum_column21_6)               //           
    );    
    
    FA FA_inst_17(
        .A              (sum_column21[0])            ,
        .B              (sum_column21[1])            ,
        .Cin            (sum_column21[2])            ,
        .sum            (sum_column21_7)            ,
        .carry          (sum_column22_5)               //           
    );    
    
    FA FA_inst_18(
        .A              (sum_column22[0])            ,
        .B              (sum_column22[1])            ,
        .Cin            (sum_column22[2])            ,
        .sum            (sum_column22_6)            ,
        .carry          (sum_column23_5)               //           
    );    
    
    FA FA_inst_19(
        .A              (sum_column23[0])            ,
        .B              (sum_column23[1])            ,
        .Cin            (sum_column23[2])            ,
        .sum            (sum_column23_6)            ,
        .carry          (sum_column24_4)               //           
    );    
    
    FA FA_inst_20(
        .A              (sum_column24[0])            ,
        .B              (sum_column24[1])            ,
        .Cin            (sum_column24[2])            ,
        .sum            (sum_column24_5)            ,
        .carry          (sum_column25_4)               //           
    );    
    
    FA FA_inst_21(
        .A              (sum_column25[0])            ,
        .B              (sum_column25[1])            ,
        .Cin            (sum_column25[2])            ,
        .sum            (sum_column25_5)            ,
        .carry          (sum_column26_3)               //           
    );    
    
    FA FA_inst_22(
        .A              (sum_column26[0])            ,
        .B              (sum_column26[1])            ,
        .Cin            (sum_column26[2])            ,
        .sum            (sum_column26_4)            ,
        .carry          (sum_column27_3)               //           
    );    
    
    FA FA_inst_23(
        .A              (sum_column27[0])            ,
        .B              (sum_column27[1])            ,
        .Cin            (sum_column27[2])            ,
        .sum            (sum_column27_4)            ,
        .carry          (sum_column28_2)               //           
    );    
    
    FA FA_inst_24(
        .A              (sum_column28[0])            ,
        .B              (sum_column28[1])            ,
        .Cin            (sum_column28_2)            ,
        .sum            (sum_column28_3)            ,
        .carry          (sum_column29_2)               //           
    );    
    
    FA FA_inst_25(
        .A              (sum_column29[0])            ,
        .B              (sum_column29[1])            ,
        .Cin            (sum_column29_2)            ,
        .sum            (sum_column29_3)            ,
        .carry          (sum_column30_1)               //           
    );    
    
    HA HA_inst_26(
        .A              (sum_column6[3])            ,
        .B              (sum_column6_4)            ,
        .sum            (sum_column6_6)            ,
        .carry          (sum_column7_6)               //           
    );   
    
    FA FA_inst_27(
        .A              (sum_column7[3])            ,
        .B              (sum_column7_4)            ,
        .Cin            (sum_column7_5)            ,
        .sum            (sum_column7_7)            ,
        .carry          (sum_column8_7)               //           
    );    
    
    FA FA_inst_28(
        .A              (sum_column8[3])            ,
        .B              (sum_column8[4])            ,
        .Cin            (sum_column8_5)            ,
        .sum            (sum_column8_8)            ,
        .carry          (sum_column9_7)               //           
    );    
    
    FA FA_inst_29(
        .A              (sum_column9[3])            ,
        .B              (sum_column9[4])            ,
        .Cin            (sum_column9_5)            ,
        .sum            (sum_column9_8)            ,
        .carry          (sum_column10_8)               //           
    );    
    
    FA FA_inst_30(
        .A              (sum_column10[3])            ,
        .B              (sum_column10[4])            ,
        .Cin            (sum_column10[5])            ,
        .sum            (sum_column10_9)            ,
        .carry          (sum_column11_8)               //           
    );    
    
    FA FA_inst_31(
        .A              (sum_column11[3])            ,
        .B              (sum_column11[4])            ,
        .Cin            (sum_column11[5])            ,
        .sum            (sum_column11_9)            ,
        .carry          (sum_column12_9)               //           
    );    
    
    FA FA_inst_32(
        .A              (sum_column12[3])            ,
        .B              (sum_column12[4])            ,
        .Cin            (sum_column12[5])            ,
        .sum            (sum_column12_10)            ,
        .carry          (sum_column13_9)               //           
    );    
    
    FA FA_inst_33(
        .A              (sum_column13[3])            ,
        .B              (sum_column13[4])            ,
        .Cin            (sum_column13[5])            ,
        .sum            (sum_column13_10)            ,
        .carry          (sum_column14_10)               //           
    );    
    
    FA FA_inst_34(
        .A              (sum_column14[3])            ,
        .B              (sum_column14[4])            ,
        .Cin            (sum_column14[5])            ,
        .sum            (sum_column14_11)            ,
        .carry          (sum_column15_10)               //           
    );    
    
    FA FA_inst_35(
        .A              (sum_column15[3])            ,
        .B              (sum_column15[4])            ,
        .Cin            (sum_column15[5])            ,
        .sum            (sum_column15_11)            ,
        .carry          (sum_column16_11)               //           
    );    
    
    FA FA_inst_36(
        .A              (sum_column16[3])            ,
        .B              (sum_column16[4])            ,
        .Cin            (sum_column16[5])            ,
        .sum            (sum_column16_12)            ,
        .carry          (sum_column17_10)               //           
    );    
    
    FA FA_inst_37(
        .A              (sum_column17[3])            ,
        .B              (sum_column17[4])            ,
        .Cin            (sum_column17[5])            ,
        .sum            (sum_column17_11)            ,
        .carry          (sum_column18_9)               //           
    );    
    
    FA FA_inst_38(
        .A              (sum_column18[3])            ,
        .B              (sum_column18[4])            ,
        .Cin            (sum_column18[5])            ,
        .sum            (sum_column18_10)            ,
        .carry          (sum_column19_9)               //           
    );    
    
    FA FA_inst_39(
        .A              (sum_column19[3])            ,
        .B              (sum_column19[4])            ,
        .Cin            (sum_column19[5])            ,
        .sum            (sum_column19_10)            ,
        .carry          (sum_column20_8)               //           
    );    
    
    FA FA_inst_40(
        .A              (sum_column20[3])            ,
        .B              (sum_column20[4])            ,
        .Cin            (sum_column20[5])            ,
        .sum            (sum_column20_9)            ,
        .carry          (sum_column21_8)               //           
    );    
    
    FA FA_inst_41(
        .A              (sum_column21[3])            ,
        .B              (sum_column21[4])            ,
        .Cin            (sum_column21[5])            ,
        .sum            (sum_column21_9)            ,
        .carry          (sum_column22_7)               //           
    );    
    
    FA FA_inst_42(
        .A              (sum_column22[3])            ,
        .B              (sum_column22[4])            ,
        .Cin            (sum_column22_5)            ,
        .sum            (sum_column22_8)            ,
        .carry          (sum_column23_7)               //           
    );    
    
    FA FA_inst_43(
        .A              (sum_column23[3])            ,
        .B              (sum_column23[4])            ,
        .Cin            (sum_column23_5)            ,
        .sum            (sum_column23_8)            ,
        .carry          (sum_column24_6)               //           
    );    
    
    FA FA_inst_44(
        .A              (sum_column24[3])            ,
        .B              (sum_column24_4)            ,
        .Cin            (sum_column24_5)            ,
        .sum            (sum_column24_7)            ,
        .carry          (sum_column25_6)               //           
    );    
    
    FA FA_inst_45(
        .A              (sum_column25[3])            ,
        .B              (sum_column25_4)            ,
        .Cin            (sum_column25_5)            ,
        .sum            (sum_column25_7)            ,
        .carry          (sum_column26_5)               //           
    );    
    
    FA FA_inst_46(
        .A              (sum_column26_3)            ,
        .B              (sum_column26_4)            ,
        .Cin            (sum_column26_5)            ,
        .sum            (sum_column26_6)            ,
        .carry          (sum_column27_5)               //           
    );    
    
    FA FA_inst_47(
        .A              (sum_column27_3)            ,
        .B              (sum_column27_4)            ,
        .Cin            (sum_column27_5)            ,
        .sum            (sum_column27_6)            ,
        .carry          (sum_column28_4)               //           
    );    
    
    HA HA_inst_48(
        .A              (sum_column8_6)            ,
        .B              (sum_column8_7)            ,
        .sum            (sum_column8_9)            ,
        .carry          (sum_column9_9)               //           
    );   
    
    FA FA_inst_49(
        .A              (sum_column9_6)            ,
        .B              (sum_column9_7)            ,
        .Cin            (sum_column9_8)            ,
        .sum            (sum_column9_10)            ,
        .carry          (sum_column10_10)               //           
    );    
    
    FA FA_inst_50(
        .A              (sum_column10_6)            ,
        .B              (sum_column10_7)            ,
        .Cin            (sum_column10_8)            ,
        .sum            (sum_column10_11)            ,
        .carry          (sum_column11_10)               //           
    );    
    
    FA FA_inst_51(
        .A              (sum_column11_6)            ,
        .B              (sum_column11_7)            ,
        .Cin            (sum_column11_8)            ,
        .sum            (sum_column11_11)            ,
        .carry          (sum_column12_11)               //           
    );    
    
    FA FA_inst_52(
        .A              (sum_column12[6])            ,
        .B              (sum_column12_7)            ,
        .Cin            (sum_column12_8)            ,
        .sum            (sum_column12_12)            ,
        .carry          (sum_column13_11)               //           
    );    
    
    FA FA_inst_53(
        .A              (sum_column13[6])            ,
        .B              (sum_column13_7)            ,
        .Cin            (sum_column13_8)            ,
        .sum            (sum_column13_12)            ,
        .carry          (sum_column14_12)               //           
    );    
    
    FA FA_inst_54(
        .A              (sum_column14[6])            ,
        .B              (sum_column14[7])            ,
        .Cin            (sum_column14_8)            ,
        .sum            (sum_column14_13)            ,
        .carry          (sum_column15_12)               //           
    );    
    
    FA FA_inst_55(
        .A              (sum_column15[6])            ,
        .B              (sum_column15[7])            ,
        .Cin            (sum_column15_8)            ,
        .sum            (sum_column15_13)            ,
        .carry          (sum_column16_13)               //           
    );    
    
    FA FA_inst_56(
        .A              (sum_column16[6])            ,
        .B              (sum_column16[7])            ,
        .Cin            (sum_column16[8])            ,
        .sum            (sum_column16_14)            ,
        .carry          (sum_column17_12)               //           
    );    
    
    FA FA_inst_57(
        .A              (sum_column17[6])            ,
        .B              (sum_column17[7])            ,
        .Cin            (sum_column17_8)            ,
        .sum            (sum_column17_13)            ,
        .carry          (sum_column18_11)               //           
    );    
    
    FA FA_inst_58(
        .A              (sum_column18[6])            ,
        .B              (sum_column18_7)            ,
        .Cin            (sum_column18_8)            ,
        .sum            (sum_column18_12)            ,
        .carry          (sum_column19_11)               //           
    );    
    
    FA FA_inst_59(
        .A              (sum_column19[6])            ,
        .B              (sum_column19_7)            ,
        .Cin            (sum_column19_8)            ,
        .sum            (sum_column19_12)            ,
        .carry          (sum_column20_10)               //           
    );    
    
    FA FA_inst_60(
        .A              (sum_column20_6)            ,
        .B              (sum_column20_7)            ,
        .Cin            (sum_column20_8)            ,
        .sum            (sum_column20_11)            ,
        .carry          (sum_column21_10)               //           
    );    
    
    FA FA_inst_61(
        .A              (sum_column21_6)            ,
        .B              (sum_column21_7)            ,
        .Cin            (sum_column21_8)            ,
        .sum            (sum_column21_11)            ,
        .carry          (sum_column22_9)               //           
    );    
    
    FA FA_inst_62(
        .A              (sum_column22_6)            ,
        .B              (sum_column22_7)            ,
        .Cin            (sum_column22_8)            ,
        .sum            (sum_column22_10)            ,
        .carry          (sum_column23_9)               //           
    );    
    
    FA FA_inst_63(
        .A              (sum_column23_6)            ,
        .B              (sum_column23_7)            ,
        .Cin            (sum_column23_8)            ,
        .sum            (sum_column23_10)            ,
        .carry          (sum_column24_8)               //           
    );    
    
    FA FA_inst_64(
        .A              (sum_column24_6)            ,
        .B              (sum_column24_7)            ,
        .Cin            (sum_column24_8)            ,
        .sum            (sum_column24_9)            ,
        .carry          (sum_column25_8)               //           
    );    
    
    FA FA_inst_65(
        .A              (sum_column25_6)            ,
        .B              (sum_column25_7)            ,
        .Cin            (sum_column25_8)            ,
        .sum            (sum_column25_9)            ,
        .carry          (sum_column26_7)               //           
    );    
    
    HA HA_inst_66(
        .A              (sum_column10_9)            ,
        .B              (sum_column10_10)            ,
        .sum            (sum_column10_12)            ,
        .carry          (sum_column11_12)               //           
    );   
    
    FA FA_inst_67(
        .A              (sum_column11_9)            ,
        .B              (sum_column11_10)            ,
        .Cin            (sum_column11_11)            ,
        .sum            (sum_column11_13)            ,
        .carry          (sum_column12_13)               //           
    );    
    
    FA FA_inst_68(
        .A              (sum_column12_9)            ,
        .B              (sum_column12_10)            ,
        .Cin            (sum_column12_11)            ,
        .sum            (sum_column12_14)            ,
        .carry          (sum_column13_13)               //           
    );    
    
    FA FA_inst_69(
        .A              (sum_column13_9)            ,
        .B              (sum_column13_10)            ,
        .Cin            (sum_column13_11)            ,
        .sum            (sum_column13_14)            ,
        .carry          (sum_column14_14)               //           
    );    
    
    FA FA_inst_70(
        .A              (sum_column14_9)            ,
        .B              (sum_column14_10)            ,
        .Cin            (sum_column14_11)            ,
        .sum            (sum_column14_15)            ,
        .carry          (sum_column15_14)               //           
    );    
    
    FA FA_inst_71(
        .A              (sum_column15_9)            ,
        .B              (sum_column15_10)            ,
        .Cin            (sum_column15_11)            ,
        .sum            (sum_column15_15)            ,
        .carry          (sum_column16_15)               //           
    );    
    
    FA FA_inst_72(
        .A              (sum_column16_9)            ,
        .B              (sum_column16_10)            ,
        .Cin            (sum_column16_11)            ,
        .sum            (sum_column16_16)            ,
        .carry          (sum_column17_14)               //           
    );    
    
    FA FA_inst_73(
        .A              (sum_column17_9)            ,
        .B              (sum_column17_10)            ,
        .Cin            (sum_column17_11)            ,
        .sum            (sum_column17_15)            ,
        .carry          (sum_column18_13)               //           
    );    
    
    FA FA_inst_74(
        .A              (sum_column18_9)            ,
        .B              (sum_column18_10)            ,
        .Cin            (sum_column18_11)            ,
        .sum            (sum_column18_14)            ,
        .carry          (sum_column19_13)               //           
    );    
    
    FA FA_inst_75(
        .A              (sum_column19_9)            ,
        .B              (sum_column19_10)            ,
        .Cin            (sum_column19_11)            ,
        .sum            (sum_column19_14)            ,
        .carry          (sum_column20_12)               //           
    );    
    
    FA FA_inst_76(
        .A              (sum_column20_9)            ,
        .B              (sum_column20_10)            ,
        .Cin            (sum_column20_11)            ,
        .sum            (sum_column20_13)            ,
        .carry          (sum_column21_12)               //           
    );    
    
    FA FA_inst_77(
        .A              (sum_column21_9)            ,
        .B              (sum_column21_10)            ,
        .Cin            (sum_column21_11)            ,
        .sum            (sum_column21_13)            ,
        .carry          (sum_column22_11)               //           
    );    
    
    FA FA_inst_78(
        .A              (sum_column22_9)            ,
        .B              (sum_column22_10)            ,
        .Cin            (sum_column22_11)            ,
        .sum            (sum_column22_12)            ,
        .carry          (sum_column23_11)               //           
    );    
    
    FA FA_inst_79(
        .A              (sum_column23_9)            ,
        .B              (sum_column23_10)            ,
        .Cin            (sum_column23_11)            ,
        .sum            (sum_column23_12)            ,
        .carry          (sum_column24_10)               //           
    );    
    
    HA HA_inst_80(
        .A              (sum_column12_12)            ,
        .B              (sum_column12_13)            ,
        .sum            (sum_column12_15)            ,
        .carry          (sum_column13_15)               //           
    );   
    
    FA FA_inst_81(
        .A              (sum_column13_12)            ,
        .B              (sum_column13_13)            ,
        .Cin            (sum_column13_14)            ,
        .sum            (sum_column13_16)            ,
        .carry          (sum_column14_16)               //           
    );    
    
    FA FA_inst_82(
        .A              (sum_column14_12)            ,
        .B              (sum_column14_13)            ,
        .Cin            (sum_column14_14)            ,
        .sum            (sum_column14_17)            ,
        .carry          (sum_column15_16)               //           
    );    
    
    FA FA_inst_83(
        .A              (sum_column15_12)            ,
        .B              (sum_column15_13)            ,
        .Cin            (sum_column15_14)            ,
        .sum            (sum_column15_17)            ,
        .carry          (sum_column16_17)               //           
    );    
    
    FA FA_inst_84(
        .A              (sum_column16_12)            ,
        .B              (sum_column16_13)            ,
        .Cin            (sum_column16_14)            ,
        .sum            (sum_column16_18)            ,
        .carry          (sum_column17_16)               //           
    );    
    
    FA FA_inst_85(
        .A              (sum_column17_12)            ,
        .B              (sum_column17_13)            ,
        .Cin            (sum_column17_14)            ,
        .sum            (sum_column17_17)            ,
        .carry          (sum_column18_15)               //           
    );    
    
    FA FA_inst_86(
        .A              (sum_column18_12)            ,
        .B              (sum_column18_13)            ,
        .Cin            (sum_column18_14)            ,
        .sum            (sum_column18_16)            ,
        .carry          (sum_column19_15)               //           
    );    
    
    FA FA_inst_87(
        .A              (sum_column19_12)            ,
        .B              (sum_column19_13)            ,
        .Cin            (sum_column19_14)            ,
        .sum            (sum_column19_16)            ,
        .carry          (sum_column20_14)               //           
    );    
    
    FA FA_inst_88(
        .A              (sum_column20_12)            ,
        .B              (sum_column20_13)            ,
        .Cin            (sum_column20_14)            ,
        .sum            (sum_column20_15)            ,
        .carry          (sum_column21_14)               //           
    );    
    
    FA FA_inst_89(
        .A              (sum_column21_12)            ,
        .B              (sum_column21_13)            ,
        .Cin            (sum_column21_14)            ,
        .sum            (sum_column21_15)            ,
        .carry          (sum_column22_13)               //           
    );    
    
    HA HA_inst_90(
        .A              (sum_column14_15)            ,
        .B              (sum_column14_16)            ,
        .sum            (sum_column14_18)            ,
        .carry          (sum_column15_18)               //           
    );   
    
    FA FA_inst_91(
        .A              (sum_column15_15)            ,
        .B              (sum_column15_16)            ,
        .Cin            (sum_column15_17)            ,
        .sum            (sum_column15_19)            ,
        .carry          (sum_column16_19)               //           
    );    
    
    FA FA_inst_92(
        .A              (sum_column16_15)            ,
        .B              (sum_column16_16)            ,
        .Cin            (sum_column16_17)            ,
        .sum            (sum_column16_20)            ,
        .carry          (sum_column17_18)               //           
    );    
    
    FA FA_inst_93(
        .A              (sum_column17_15)            ,
        .B              (sum_column17_16)            ,
        .Cin            (sum_column17_17)            ,
        .sum            (sum_column17_19)            ,
        .carry          (sum_column18_17)               //           
    );    
    
    FA FA_inst_94(
        .A              (sum_column18_15)            ,
        .B              (sum_column18_16)            ,
        .Cin            (sum_column18_17)            ,
        .sum            (sum_column18_18)            ,
        .carry          (sum_column19_17)               //           
    );    
    
    FA FA_inst_95(
        .A              (sum_column19_15)            ,
        .B              (sum_column19_16)            ,
        .Cin            (sum_column19_17)            ,
        .sum            (sum_column19_18)            ,
        .carry          (sum_column20_16)               //           
    );    
    
    HA HA_inst_96(
        .A              (sum_column16_18)            ,
        .B              (sum_column16_19)            ,
        .sum            (sum_column16_21)            ,
        .carry          (sum_column17_20)               //           
    );   
    
    FA FA_inst_97(
        .A              (sum_column17_18)            ,
        .B              (sum_column17_19)            ,
        .Cin            (sum_column17_20)            ,
        .sum            (sum_column17_21)            ,
        .carry          (sum_column18_19)               //           
    );    
    

	assign vector0 = {
        sum_column31[0]				,				
		sum_column30[0]				,				
		1'b0							,				
		sum_column28_3				,				
		1'b0							,				
		sum_column26_6				,				
		1'b0							,				
		sum_column24_9				,				
		1'b0							,				
		sum_column22_12				,				
		1'b0							,				
		sum_column20_15				,				
		1'b0							,				
		sum_column18_18				,				
		1'b0							,				
		sum_column16_20				,				
		sum_column15_18				,				
		sum_column14_17				,				
		sum_column13_15				,				
		sum_column12_14				,				
		sum_column11_12				,				
		sum_column10_11				,				
		sum_column9_9				,				
		sum_column8_8				,				
		sum_column7_6				,				
		sum_column6_5				,				
		sum_column5_3				,				
		sum_column4[2]				,				
		sum_column3[0]				,				
		sum_column2[0]				,				
		sum_column1[0]				,				
		sum_column0[0]								

    };
    assign vector1 = {
        sum_column31[1]				,				
		sum_column30_1				,				
		sum_column29_3				,				
		sum_column28_4				,				
		sum_column27_6				,				
		sum_column26_7				,				
		sum_column25_9				,				
		sum_column24_10				,				
		sum_column23_12				,				
		sum_column22_13				,				
		sum_column21_15				,				
		sum_column20_16				,				
		sum_column19_18				,				
		sum_column18_19				,				
		sum_column17_21				,				
		sum_column16_21				,				
		sum_column15_19				,				
		sum_column14_18				,				
		sum_column13_16				,				
		sum_column12_15				,				
		sum_column11_13				,				
		sum_column10_12				,				
		sum_column9_10				,				
		sum_column8_9				,				
		sum_column7_7				,				
		sum_column6_6				,				
		sum_column5_4				,				
		sum_column4_3				,				
		sum_column3[1]				,				
		sum_column2[1]				,				
		1'b0						,				
		1'b0										

    };

    

endmodule

