`timescale 1ns/1ns
module adder<#width1>(
    input           [<#width1>:1]      A                 ,
    input           [<#width1>:1]      B                 ,
    input                       c0                ,
    output          [<#width1>:1]      S                 ,
    output                      c<#width1>               
);

    <wire definition>

    <adder4 instantiation>


endmodule

